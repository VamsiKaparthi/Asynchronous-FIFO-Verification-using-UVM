package pkg;
        `include "uvm_macros.svh"
        import uvm_pkg::*;
        `include "define.svh"
        `include "seq_item.sv"
        `include "sequencer.sv"
        `include "sequence.sv"
  `include "wr_driver.sv"
        `include "rd_driver.sv"
        `include "wr_monitor.sv"
        `include "rd_monitor.sv"
        `include "write_agent.sv"
        `include "read_agent.sv"
        `include "scoreboard.sv"
        `include "coverage.sv"
        `include "environment.sv"
        `include "test.sv"
endpackage
