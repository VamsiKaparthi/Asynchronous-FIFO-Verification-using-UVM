parameter DSIZE = 8;
parameter ASIZE = 4;
parameter DEPTH = 1<<ASIZE;
parameter N = 100;
